package shared_pkg;
	typedef enum logic {SHIFT, ROTATE} mode_e;
	typedef enum logic {RIGHT, LEFT} direction_e;
endpackage : shared_pkg